

module weights_luts #(N1=98, N2=10, W_K=4)(
  output wire [W_K-1:0] weights_n1_mag [N1/2][N2],
  output wire [W_K-1:0] weights_n1_pol [N1/2][N2],
  output wire [W_K-1:0] weights_n2 [N2]
);
  assign weights_n1_mag = '{
    '{ 4'd12     , 4'd15     , 4'd5      , 4'd0      , 4'd3      , 4'd11     , 4'd3      , 4'd7      , 4'd9      , 4'd3       },
    '{ 4'd5      , 4'd2      , 4'd4      , 4'd7      , 4'd6      , 4'd8      , 4'd8      , 4'd12     , 4'd10     , 4'd1       },
    '{ 4'd6      , 4'd7      , 4'd7      , 4'd14     , 4'd8      , 4'd1      , 4'd5      , 4'd9      , 4'd13     , 4'd8       },
    '{ 4'd9      , 4'd4      , 4'd3      , 4'd0      , 4'd3      , 4'd5      , 4'd14     , 4'd15     , 4'd15     , 4'd0       },
    '{ 4'd2      , 4'd3      , 4'd8      , 4'd1      , 4'd3      , 4'd13     , 4'd3      , 4'd3      , 4'd14     , 4'd7       },
    '{ 4'd0      , 4'd1      , 4'd9      , 4'd9      , 4'd15     , 4'd0      , 4'd15     , 4'd10     , 4'd4      , 4'd7       },
    '{ 4'd3      , 4'd14     , 4'd11     , 4'd2      , 4'd7      , 4'd12     , 4'd2      , 4'd0      , 4'd0      , 4'd4       },
    '{ 4'd5      , 4'd5      , 4'd6      , 4'd8      , 4'd4      , 4'd1      , 4'd15     , 4'd4      , 4'd9      , 4'd10      },
    '{ 4'd10     , 4'd15     , 4'd8      , 4'd1      , 4'd1      , 4'd7      , 4'd9      , 4'd9      , 4'd3      , 4'd6       },
    '{ 4'd7      , 4'd11     , 4'd14     , 4'd2      , 4'd11     , 4'd0      , 4'd14     , 4'd3      , 4'd5      , 4'd12      },
    '{ 4'd9      , 4'd10     , 4'd4      , 4'd11     , 4'd4      , 4'd6      , 4'd4      , 4'd15     , 4'd15     , 4'd4       },
    '{ 4'd3      , 4'd12     , 4'd4      , 4'd4      , 4'd8      , 4'd14     , 4'd15     , 4'd4      , 4'd3      , 4'd10      },
    '{ 4'd7      , 4'd15     , 4'd13     , 4'd5      , 4'd5      , 4'd0      , 4'd1      , 4'd5      , 4'd9      , 4'd3       },
    '{ 4'd0      , 4'd15     , 4'd5      , 4'd14     , 4'd0      , 4'd1      , 4'd2      , 4'd4      , 4'd2      , 4'd0       },
    '{ 4'd13     , 4'd3      , 4'd2      , 4'd10     , 4'd13     , 4'd0      , 4'd7      , 4'd5      , 4'd9      , 4'd15      },
    '{ 4'd0      , 4'd10     , 4'd2      , 4'd11     , 4'd10     , 4'd15     , 4'd7      , 4'd11     , 4'd2      , 4'd9       },
    '{ 4'd2      , 4'd14     , 4'd3      , 4'd14     , 4'd11     , 4'd3      , 4'd2      , 4'd14     , 4'd3      , 4'd4       },
    '{ 4'd1      , 4'd2      , 4'd11     , 4'd14     , 4'd9      , 4'd10     , 4'd1      , 4'd4      , 4'd10     , 4'd6       },
    '{ 4'd11     , 4'd8      , 4'd11     , 4'd2      , 4'd3      , 4'd0      , 4'd0      , 4'd6      , 4'd0      , 4'd6       },
    '{ 4'd3      , 4'd14     , 4'd10     , 4'd3      , 4'd8      , 4'd12     , 4'd8      , 4'd13     , 4'd14     , 4'd8       },
    '{ 4'd13     , 4'd2      , 4'd3      , 4'd14     , 4'd2      , 4'd11     , 4'd13     , 4'd0      , 4'd8      , 4'd8       },
    '{ 4'd3      , 4'd15     , 4'd8      , 4'd10     , 4'd2      , 4'd8      , 4'd4      , 4'd3      , 4'd12     , 4'd13      },
    '{ 4'd14     , 4'd0      , 4'd4      , 4'd3      , 4'd13     , 4'd11     , 4'd12     , 4'd6      , 4'd13     , 4'd9       },
    '{ 4'd13     , 4'd11     , 4'd8      , 4'd0      , 4'd8      , 4'd13     , 4'd5      , 4'd14     , 4'd9      , 4'd0       },
    '{ 4'd12     , 4'd9      , 4'd6      , 4'd5      , 4'd13     , 4'd3      , 4'd1      , 4'd8      , 4'd0      , 4'd4       },
    '{ 4'd11     , 4'd11     , 4'd9      , 4'd6      , 4'd5      , 4'd15     , 4'd13     , 4'd7      , 4'd8      , 4'd8       },
    '{ 4'd15     , 4'd9      , 4'd2      , 4'd8      , 4'd6      , 4'd15     , 4'd11     , 4'd6      , 4'd15     , 4'd13      },
    '{ 4'd9      , 4'd1      , 4'd15     , 4'd6      , 4'd12     , 4'd8      , 4'd13     , 4'd8      , 4'd3      , 4'd2       },
    '{ 4'd15     , 4'd3      , 4'd10     , 4'd12     , 4'd6      , 4'd3      , 4'd6      , 4'd14     , 4'd13     , 4'd5       },
    '{ 4'd7      , 4'd11     , 4'd0      , 4'd11     , 4'd8      , 4'd4      , 4'd10     , 4'd6      , 4'd11     , 4'd5       },
    '{ 4'd13     , 4'd12     , 4'd15     , 4'd8      , 4'd2      , 4'd11     , 4'd3      , 4'd9      , 4'd7      , 4'd5       },
    '{ 4'd3      , 4'd14     , 4'd4      , 4'd5      , 4'd13     , 4'd3      , 4'd3      , 4'd7      , 4'd9      , 4'd9       },
    '{ 4'd9      , 4'd7      , 4'd3      , 4'd14     , 4'd10     , 4'd2      , 4'd12     , 4'd3      , 4'd15     , 4'd9       },
    '{ 4'd10     , 4'd11     , 4'd13     , 4'd7      , 4'd7      , 4'd13     , 4'd5      , 4'd1      , 4'd12     , 4'd2       },
    '{ 4'd2      , 4'd8      , 4'd1      , 4'd5      , 4'd8      , 4'd15     , 4'd4      , 4'd0      , 4'd11     , 4'd2       },
    '{ 4'd5      , 4'd14     , 4'd5      , 4'd14     , 4'd0      , 4'd14     , 4'd8      , 4'd13     , 4'd1      , 4'd1       },
    '{ 4'd0      , 4'd3      , 4'd8      , 4'd11     , 4'd8      , 4'd4      , 4'd4      , 4'd0      , 4'd9      , 4'd3       },
    '{ 4'd7      , 4'd12     , 4'd3      , 4'd2      , 4'd14     , 4'd13     , 4'd1      , 4'd1      , 4'd2      , 4'd1       },
    '{ 4'd13     , 4'd4      , 4'd13     , 4'd2      , 4'd5      , 4'd5      , 4'd12     , 4'd12     , 4'd5      , 4'd13      },
    '{ 4'd2      , 4'd15     , 4'd11     , 4'd5      , 4'd7      , 4'd7      , 4'd11     , 4'd6      , 4'd14     , 4'd1       },
    '{ 4'd6      , 4'd7      , 4'd2      , 4'd12     , 4'd11     , 4'd3      , 4'd1      , 4'd9      , 4'd13     , 4'd14      },
    '{ 4'd5      , 4'd9      , 4'd9      , 4'd2      , 4'd0      , 4'd11     , 4'd9      , 4'd12     , 4'd11     , 4'd1       },
    '{ 4'd9      , 4'd10     , 4'd0      , 4'd6      , 4'd15     , 4'd0      , 4'd10     , 4'd4      , 4'd14     , 4'd8       },
    '{ 4'd4      , 4'd15     , 4'd3      , 4'd3      , 4'd8      , 4'd8      , 4'd11     , 4'd13     , 4'd11     , 4'd14      },
    '{ 4'd7      , 4'd0      , 4'd3      , 4'd8      , 4'd7      , 4'd7      , 4'd13     , 4'd10     , 4'd1      , 4'd8       },
    '{ 4'd4      , 4'd7      , 4'd0      , 4'd11     , 4'd12     , 4'd4      , 4'd9      , 4'd0      , 4'd10     , 4'd14      },
    '{ 4'd6      , 4'd12     , 4'd4      , 4'd2      , 4'd4      , 4'd6      , 4'd3      , 4'd10     , 4'd3      , 4'd7       },
    '{ 4'd8      , 4'd13     , 4'd13     , 4'd5      , 4'd0      , 4'd8      , 4'd15     , 4'd15     , 4'd5      , 4'd11      },
    '{ 4'd4      , 4'd7      , 4'd12     , 4'd13     , 4'd10     , 4'd10     , 4'd4      , 4'd14     , 4'd1      , 4'd11      }
  };

  assign weights_n1_pol = '{
    '{ 4'd3      , 4'd3      , 4'd9      , 4'd2      , 4'd5      , 4'd2      , 4'd3      , 4'd14     , 4'd5      , 4'd10      },
    '{ 4'd11     , 4'd7      , 4'd12     , 4'd12     , 4'd2      , 4'd13     , 4'd7      , 4'd1      , 4'd6      , 4'd10      },
    '{ 4'd5      , 4'd0      , 4'd14     , 4'd11     , 4'd0      , 4'd10     , 4'd12     , 4'd3      , 4'd10     , 4'd1       },
    '{ 4'd10     , 4'd9      , 4'd12     , 4'd13     , 4'd9      , 4'd6      , 4'd6      , 4'd7      , 4'd8      , 4'd13      },
    '{ 4'd8      , 4'd7      , 4'd0      , 4'd8      , 4'd6      , 4'd8      , 4'd15     , 4'd9      , 4'd8      , 4'd3       },
    '{ 4'd6      , 4'd1      , 4'd7      , 4'd4      , 4'd9      , 4'd2      , 4'd12     , 4'd0      , 4'd8      , 4'd2       },
    '{ 4'd13     , 4'd7      , 4'd8      , 4'd4      , 4'd4      , 4'd12     , 4'd1      , 4'd7      , 4'd14     , 4'd6       },
    '{ 4'd9      , 4'd4      , 4'd1      , 4'd5      , 4'd9      , 4'd7      , 4'd11     , 4'd13     , 4'd1      , 4'd3       },
    '{ 4'd5      , 4'd7      , 4'd3      , 4'd6      , 4'd6      , 4'd7      , 4'd9      , 4'd1      , 4'd9      , 4'd6       },
    '{ 4'd0      , 4'd3      , 4'd8      , 4'd4      , 4'd1      , 4'd4      , 4'd5      , 4'd0      , 4'd3      , 4'd14      },
    '{ 4'd10     , 4'd1      , 4'd4      , 4'd4      , 4'd4      , 4'd0      , 4'd0      , 4'd15     , 4'd10     , 4'd13      },
    '{ 4'd8      , 4'd14     , 4'd11     , 4'd11     , 4'd15     , 4'd15     , 4'd4      , 4'd6      , 4'd9      , 4'd12      },
    '{ 4'd11     , 4'd15     , 4'd3      , 4'd3      , 4'd12     , 4'd2      , 4'd1      , 4'd10     , 4'd2      , 4'd1       },
    '{ 4'd11     , 4'd3      , 4'd12     , 4'd4      , 4'd10     , 4'd1      , 4'd1      , 4'd0      , 4'd7      , 4'd8       },
    '{ 4'd10     , 4'd4      , 4'd3      , 4'd5      , 4'd6      , 4'd3      , 4'd2      , 4'd9      , 4'd8      , 4'd12      },
    '{ 4'd1      , 4'd12     , 4'd4      , 4'd10     , 4'd0      , 4'd8      , 4'd13     , 4'd3      , 4'd9      , 4'd5       },
    '{ 4'd5      , 4'd1      , 4'd7      , 4'd13     , 4'd14     , 4'd8      , 4'd6      , 4'd4      , 4'd7      , 4'd3       },
    '{ 4'd5      , 4'd11     , 4'd12     , 4'd3      , 4'd6      , 4'd4      , 4'd7      , 4'd3      , 4'd15     , 4'd0       },
    '{ 4'd5      , 4'd11     , 4'd11     , 4'd14     , 4'd9      , 4'd3      , 4'd7      , 4'd5      , 4'd5      , 4'd12      },
    '{ 4'd8      , 4'd11     , 4'd14     , 4'd0      , 4'd8      , 4'd3      , 4'd6      , 4'd9      , 4'd10     , 4'd3       },
    '{ 4'd2      , 4'd11     , 4'd7      , 4'd0      , 4'd3      , 4'd10     , 4'd14     , 4'd0      , 4'd3      , 4'd6       },
    '{ 4'd1      , 4'd12     , 4'd11     , 4'd9      , 4'd2      , 4'd13     , 4'd9      , 4'd4      , 4'd9      , 4'd13      },
    '{ 4'd11     , 4'd1      , 4'd3      , 4'd2      , 4'd4      , 4'd13     , 4'd9      , 4'd15     , 4'd7      , 4'd4       },
    '{ 4'd9      , 4'd14     , 4'd4      , 4'd1      , 4'd2      , 4'd13     , 4'd14     , 4'd13     , 4'd7      , 4'd2       },
    '{ 4'd3      , 4'd9      , 4'd10     , 4'd7      , 4'd10     , 4'd6      , 4'd6      , 4'd12     , 4'd15     , 4'd2       },
    '{ 4'd10     , 4'd3      , 4'd6      , 4'd14     , 4'd0      , 4'd13     , 4'd12     , 4'd15     , 4'd10     , 4'd8       },
    '{ 4'd0      , 4'd10     , 4'd11     , 4'd13     , 4'd7      , 4'd14     , 4'd6      , 4'd13     , 4'd5      , 4'd14      },
    '{ 4'd15     , 4'd9      , 4'd6      , 4'd5      , 4'd11     , 4'd2      , 4'd7      , 4'd12     , 4'd1      , 4'd9       },
    '{ 4'd2      , 4'd2      , 4'd12     , 4'd14     , 4'd5      , 4'd11     , 4'd6      , 4'd4      , 4'd15     , 4'd13      },
    '{ 4'd2      , 4'd12     , 4'd14     , 4'd13     , 4'd2      , 4'd1      , 4'd12     , 4'd0      , 4'd9      , 4'd0       },
    '{ 4'd2      , 4'd8      , 4'd3      , 4'd13     , 4'd10     , 4'd0      , 4'd10     , 4'd11     , 4'd8      , 4'd8       },
    '{ 4'd1      , 4'd0      , 4'd5      , 4'd8      , 4'd2      , 4'd15     , 4'd3      , 4'd12     , 4'd14     , 4'd5       },
    '{ 4'd11     , 4'd3      , 4'd8      , 4'd6      , 4'd4      , 4'd6      , 4'd12     , 4'd3      , 4'd6      , 4'd2       },
    '{ 4'd12     , 4'd12     , 4'd6      , 4'd5      , 4'd11     , 4'd5      , 4'd13     , 4'd9      , 4'd4      , 4'd6       },
    '{ 4'd13     , 4'd5      , 4'd11     , 4'd15     , 4'd1      , 4'd3      , 4'd13     , 4'd3      , 4'd10     , 4'd8       },
    '{ 4'd14     , 4'd9      , 4'd5      , 4'd13     , 4'd5      , 4'd6      , 4'd0      , 4'd9      , 4'd14     , 4'd7       },
    '{ 4'd5      , 4'd15     , 4'd1      , 4'd5      , 4'd6      , 4'd12     , 4'd10     , 4'd10     , 4'd11     , 4'd6       },
    '{ 4'd14     , 4'd14     , 4'd8      , 4'd7      , 4'd13     , 4'd5      , 4'd15     , 4'd11     , 4'd10     , 4'd3       },
    '{ 4'd10     , 4'd2      , 4'd9      , 4'd11     , 4'd9      , 4'd3      , 4'd13     , 4'd14     , 4'd2      , 4'd5       },
    '{ 4'd10     , 4'd4      , 4'd1      , 4'd5      , 4'd15     , 4'd14     , 4'd8      , 4'd3      , 4'd5      , 4'd8       },
    '{ 4'd4      , 4'd10     , 4'd1      , 4'd7      , 4'd8      , 4'd1      , 4'd2      , 4'd1      , 4'd14     , 4'd1       },
    '{ 4'd7      , 4'd5      , 4'd11     , 4'd14     , 4'd0      , 4'd4      , 4'd15     , 4'd1      , 4'd1      , 4'd13      },
    '{ 4'd12     , 4'd6      , 4'd14     , 4'd6      , 4'd0      , 4'd2      , 4'd3      , 4'd7      , 4'd12     , 4'd9       },
    '{ 4'd14     , 4'd2      , 4'd11     , 4'd4      , 4'd9      , 4'd14     , 4'd0      , 4'd12     , 4'd6      , 4'd9       },
    '{ 4'd2      , 4'd4      , 4'd7      , 4'd3      , 4'd0      , 4'd12     , 4'd5      , 4'd4      , 4'd13     , 4'd0       },
    '{ 4'd13     , 4'd2      , 4'd3      , 4'd1      , 4'd7      , 4'd10     , 4'd1      , 4'd14     , 4'd13     , 4'd3       },
    '{ 4'd10     , 4'd4      , 4'd10     , 4'd1      , 4'd7      , 4'd4      , 4'd0      , 4'd10     , 4'd2      , 4'd12      },
    '{ 4'd10     , 4'd7      , 4'd4      , 4'd0      , 4'd2      , 4'd6      , 4'd9      , 4'd2      , 4'd4      , 4'd12      },
    '{ 4'd9      , 4'd9      , 4'd12     , 4'd5      , 4'd4      , 4'd10     , 4'd4      , 4'd9      , 4'd10     , 4'd12      }
  };

  assign weights_n2 = '{
    4'd9 ,
    4'd9 ,
    4'd12,
    4'd5 ,
    4'd4 ,
    4'd10,
    4'd4 ,
    4'd9 ,
    4'd10,
    4'd12
  };
endmodule
