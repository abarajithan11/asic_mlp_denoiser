
`timescale 1ns/1ps

module luts #(N1=98, N2=10, W_K=4, W_OUT=16)(
  output wire [N2-1:0][N1/2:0][W_K-1:0] weights_n1_mag,
  output wire [N2-1:0][N1/2:0][W_K-1:0] weights_n1_pol,
  output wire [N2  :0][W_K-1:0] weights_n2,
  output wire [2**W_K-1:0][W_OUT-1:0] tanh 
);
  assign weights_n1_mag = '{
    '{ 4'd12     , 4'd15     , 4'd5      , 4'd0      , 4'd3      , 4'd11     , 4'd3      , 4'd7      , 4'd9      , 4'd3      , 4'd5      , 4'd2      , 4'd4      , 4'd7      , 4'd6      , 4'd8      , 4'd8      , 4'd12     , 4'd10     , 4'd1      , 4'd6      , 4'd7      , 4'd7      , 4'd14     , 4'd8      , 4'd1      , 4'd5      , 4'd9      , 4'd13     , 4'd8      , 4'd9      , 4'd4      , 4'd3      , 4'd0      , 4'd3      , 4'd5      , 4'd14     , 4'd15     , 4'd15     , 4'd0      , 4'd2      , 4'd3      , 4'd8      , 4'd1      , 4'd3      , 4'd13     , 4'd3      , 4'd3      , 4'd14     , 4'd7       },
    '{ 4'd0      , 4'd1      , 4'd9      , 4'd9      , 4'd15     , 4'd0      , 4'd15     , 4'd10     , 4'd4      , 4'd7      , 4'd3      , 4'd14     , 4'd11     , 4'd2      , 4'd7      , 4'd12     , 4'd2      , 4'd0      , 4'd0      , 4'd4      , 4'd5      , 4'd5      , 4'd6      , 4'd8      , 4'd4      , 4'd1      , 4'd15     , 4'd4      , 4'd9      , 4'd10     , 4'd10     , 4'd15     , 4'd8      , 4'd1      , 4'd1      , 4'd7      , 4'd9      , 4'd9      , 4'd3      , 4'd6      , 4'd7      , 4'd11     , 4'd14     , 4'd2      , 4'd11     , 4'd0      , 4'd14     , 4'd3      , 4'd5      , 4'd12      },
    '{ 4'd9      , 4'd10     , 4'd4      , 4'd11     , 4'd4      , 4'd6      , 4'd4      , 4'd15     , 4'd15     , 4'd4      , 4'd3      , 4'd12     , 4'd4      , 4'd4      , 4'd8      , 4'd14     , 4'd15     , 4'd4      , 4'd3      , 4'd10     , 4'd7      , 4'd15     , 4'd13     , 4'd5      , 4'd5      , 4'd0      , 4'd1      , 4'd5      , 4'd9      , 4'd3      , 4'd0      , 4'd15     , 4'd5      , 4'd14     , 4'd0      , 4'd1      , 4'd2      , 4'd4      , 4'd2      , 4'd0      , 4'd13     , 4'd3      , 4'd2      , 4'd10     , 4'd13     , 4'd0      , 4'd7      , 4'd5      , 4'd9      , 4'd15      },
    '{ 4'd0      , 4'd10     , 4'd2      , 4'd11     , 4'd10     , 4'd15     , 4'd7      , 4'd11     , 4'd2      , 4'd9      , 4'd2      , 4'd14     , 4'd3      , 4'd14     , 4'd11     , 4'd3      , 4'd2      , 4'd14     , 4'd3      , 4'd4      , 4'd1      , 4'd2      , 4'd11     , 4'd14     , 4'd9      , 4'd10     , 4'd1      , 4'd4      , 4'd10     , 4'd6      , 4'd11     , 4'd8      , 4'd11     , 4'd2      , 4'd3      , 4'd0      , 4'd0      , 4'd6      , 4'd0      , 4'd6      , 4'd3      , 4'd14     , 4'd10     , 4'd3      , 4'd8      , 4'd12     , 4'd8      , 4'd13     , 4'd14     , 4'd8       },
    '{ 4'd13     , 4'd2      , 4'd3      , 4'd14     , 4'd2      , 4'd11     , 4'd13     , 4'd0      , 4'd8      , 4'd8      , 4'd3      , 4'd15     , 4'd8      , 4'd10     , 4'd2      , 4'd8      , 4'd4      , 4'd3      , 4'd12     , 4'd13     , 4'd14     , 4'd0      , 4'd4      , 4'd3      , 4'd13     , 4'd11     , 4'd12     , 4'd6      , 4'd13     , 4'd9      , 4'd13     , 4'd11     , 4'd8      , 4'd0      , 4'd8      , 4'd13     , 4'd5      , 4'd14     , 4'd9      , 4'd0      , 4'd12     , 4'd9      , 4'd6      , 4'd5      , 4'd13     , 4'd3      , 4'd1      , 4'd8      , 4'd0      , 4'd4       },
    '{ 4'd11     , 4'd11     , 4'd9      , 4'd6      , 4'd5      , 4'd15     , 4'd13     , 4'd7      , 4'd8      , 4'd8      , 4'd15     , 4'd9      , 4'd2      , 4'd8      , 4'd6      , 4'd15     , 4'd11     , 4'd6      , 4'd15     , 4'd13     , 4'd9      , 4'd1      , 4'd15     , 4'd6      , 4'd12     , 4'd8      , 4'd13     , 4'd8      , 4'd3      , 4'd2      , 4'd15     , 4'd3      , 4'd10     , 4'd12     , 4'd6      , 4'd3      , 4'd6      , 4'd14     , 4'd13     , 4'd5      , 4'd7      , 4'd11     , 4'd0      , 4'd11     , 4'd8      , 4'd4      , 4'd10     , 4'd6      , 4'd11     , 4'd5       },
    '{ 4'd13     , 4'd12     , 4'd15     , 4'd8      , 4'd2      , 4'd11     , 4'd3      , 4'd9      , 4'd7      , 4'd5      , 4'd3      , 4'd14     , 4'd4      , 4'd5      , 4'd13     , 4'd3      , 4'd3      , 4'd7      , 4'd9      , 4'd9      , 4'd9      , 4'd7      , 4'd3      , 4'd14     , 4'd10     , 4'd2      , 4'd12     , 4'd3      , 4'd15     , 4'd9      , 4'd10     , 4'd11     , 4'd13     , 4'd7      , 4'd7      , 4'd13     , 4'd5      , 4'd1      , 4'd12     , 4'd2      , 4'd2      , 4'd8      , 4'd1      , 4'd5      , 4'd8      , 4'd15     , 4'd4      , 4'd0      , 4'd11     , 4'd2       },
    '{ 4'd5      , 4'd14     , 4'd5      , 4'd14     , 4'd0      , 4'd14     , 4'd8      , 4'd13     , 4'd1      , 4'd1      , 4'd0      , 4'd3      , 4'd8      , 4'd11     , 4'd8      , 4'd4      , 4'd4      , 4'd0      , 4'd9      , 4'd3      , 4'd7      , 4'd12     , 4'd3      , 4'd2      , 4'd14     , 4'd13     , 4'd1      , 4'd1      , 4'd2      , 4'd1      , 4'd13     , 4'd4      , 4'd13     , 4'd2      , 4'd5      , 4'd5      , 4'd12     , 4'd12     , 4'd5      , 4'd13     , 4'd2      , 4'd15     , 4'd11     , 4'd5      , 4'd7      , 4'd7      , 4'd11     , 4'd6      , 4'd14     , 4'd1       },
    '{ 4'd6      , 4'd7      , 4'd2      , 4'd12     , 4'd11     , 4'd3      , 4'd1      , 4'd9      , 4'd13     , 4'd14     , 4'd5      , 4'd9      , 4'd9      , 4'd2      , 4'd0      , 4'd11     , 4'd9      , 4'd12     , 4'd11     , 4'd1      , 4'd9      , 4'd10     , 4'd0      , 4'd6      , 4'd15     , 4'd0      , 4'd10     , 4'd4      , 4'd14     , 4'd8      , 4'd4      , 4'd15     , 4'd3      , 4'd3      , 4'd8      , 4'd8      , 4'd11     , 4'd13     , 4'd11     , 4'd14     , 4'd7      , 4'd0      , 4'd3      , 4'd8      , 4'd7      , 4'd7      , 4'd13     , 4'd10     , 4'd1      , 4'd8       },
    '{ 4'd4      , 4'd7      , 4'd0      , 4'd11     , 4'd12     , 4'd4      , 4'd9      , 4'd0      , 4'd10     , 4'd14     , 4'd6      , 4'd12     , 4'd4      , 4'd2      , 4'd4      , 4'd6      , 4'd3      , 4'd10     , 4'd3      , 4'd7      , 4'd8      , 4'd13     , 4'd13     , 4'd5      , 4'd0      , 4'd8      , 4'd15     , 4'd15     , 4'd5      , 4'd11     , 4'd4      , 4'd7      , 4'd12     , 4'd13     , 4'd10     , 4'd10     , 4'd4      , 4'd14     , 4'd1      , 4'd11     , 4'd3      , 4'd3      , 4'd9      , 4'd2      , 4'd5      , 4'd2      , 4'd3      , 4'd14     , 4'd5      , 4'd10      }
  };

  assign weights_n1_pol = '{
    '{ 4'd11     , 4'd7      , 4'd12     , 4'd12     , 4'd2      , 4'd13     , 4'd7      , 4'd1      , 4'd6      , 4'd10     , 4'd5      , 4'd0      , 4'd14     , 4'd11     , 4'd0      , 4'd10     , 4'd12     , 4'd3      , 4'd10     , 4'd1      , 4'd10     , 4'd9      , 4'd12     , 4'd13     , 4'd9      , 4'd6      , 4'd6      , 4'd7      , 4'd8      , 4'd13     , 4'd8      , 4'd7      , 4'd0      , 4'd8      , 4'd6      , 4'd8      , 4'd15     , 4'd9      , 4'd8      , 4'd3      , 4'd6      , 4'd1      , 4'd7      , 4'd4      , 4'd9      , 4'd2      , 4'd12     , 4'd0      , 4'd8      , 4'd2       },
    '{ 4'd13     , 4'd7      , 4'd8      , 4'd4      , 4'd4      , 4'd12     , 4'd1      , 4'd7      , 4'd14     , 4'd6      , 4'd9      , 4'd4      , 4'd1      , 4'd5      , 4'd9      , 4'd7      , 4'd11     , 4'd13     , 4'd1      , 4'd3      , 4'd5      , 4'd7      , 4'd3      , 4'd6      , 4'd6      , 4'd7      , 4'd9      , 4'd1      , 4'd9      , 4'd6      , 4'd0      , 4'd3      , 4'd8      , 4'd4      , 4'd1      , 4'd4      , 4'd5      , 4'd0      , 4'd3      , 4'd14     , 4'd10     , 4'd1      , 4'd4      , 4'd4      , 4'd4      , 4'd0      , 4'd0      , 4'd15     , 4'd10     , 4'd13      },
    '{ 4'd8      , 4'd14     , 4'd11     , 4'd11     , 4'd15     , 4'd15     , 4'd4      , 4'd6      , 4'd9      , 4'd12     , 4'd11     , 4'd15     , 4'd3      , 4'd3      , 4'd12     , 4'd2      , 4'd1      , 4'd10     , 4'd2      , 4'd1      , 4'd11     , 4'd3      , 4'd12     , 4'd4      , 4'd10     , 4'd1      , 4'd1      , 4'd0      , 4'd7      , 4'd8      , 4'd10     , 4'd4      , 4'd3      , 4'd5      , 4'd6      , 4'd3      , 4'd2      , 4'd9      , 4'd8      , 4'd12     , 4'd1      , 4'd12     , 4'd4      , 4'd10     , 4'd0      , 4'd8      , 4'd13     , 4'd3      , 4'd9      , 4'd5       },
    '{ 4'd5      , 4'd1      , 4'd7      , 4'd13     , 4'd14     , 4'd8      , 4'd6      , 4'd4      , 4'd7      , 4'd3      , 4'd5      , 4'd11     , 4'd12     , 4'd3      , 4'd6      , 4'd4      , 4'd7      , 4'd3      , 4'd15     , 4'd0      , 4'd5      , 4'd11     , 4'd11     , 4'd14     , 4'd9      , 4'd3      , 4'd7      , 4'd5      , 4'd5      , 4'd12     , 4'd8      , 4'd11     , 4'd14     , 4'd0      , 4'd8      , 4'd3      , 4'd6      , 4'd9      , 4'd10     , 4'd3      , 4'd2      , 4'd11     , 4'd7      , 4'd0      , 4'd3      , 4'd10     , 4'd14     , 4'd0      , 4'd3      , 4'd6       },
    '{ 4'd1      , 4'd12     , 4'd11     , 4'd9      , 4'd2      , 4'd13     , 4'd9      , 4'd4      , 4'd9      , 4'd13     , 4'd11     , 4'd1      , 4'd3      , 4'd2      , 4'd4      , 4'd13     , 4'd9      , 4'd15     , 4'd7      , 4'd4      , 4'd9      , 4'd14     , 4'd4      , 4'd1      , 4'd2      , 4'd13     , 4'd14     , 4'd13     , 4'd7      , 4'd2      , 4'd3      , 4'd9      , 4'd10     , 4'd7      , 4'd10     , 4'd6      , 4'd6      , 4'd12     , 4'd15     , 4'd2      , 4'd10     , 4'd3      , 4'd6      , 4'd14     , 4'd0      , 4'd13     , 4'd12     , 4'd15     , 4'd10     , 4'd8       },
    '{ 4'd0      , 4'd10     , 4'd11     , 4'd13     , 4'd7      , 4'd14     , 4'd6      , 4'd13     , 4'd5      , 4'd14     , 4'd15     , 4'd9      , 4'd6      , 4'd5      , 4'd11     , 4'd2      , 4'd7      , 4'd12     , 4'd1      , 4'd9      , 4'd2      , 4'd2      , 4'd12     , 4'd14     , 4'd5      , 4'd11     , 4'd6      , 4'd4      , 4'd15     , 4'd13     , 4'd2      , 4'd12     , 4'd14     , 4'd13     , 4'd2      , 4'd1      , 4'd12     , 4'd0      , 4'd9      , 4'd0      , 4'd2      , 4'd8      , 4'd3      , 4'd13     , 4'd10     , 4'd0      , 4'd10     , 4'd11     , 4'd8      , 4'd8       },
    '{ 4'd1      , 4'd0      , 4'd5      , 4'd8      , 4'd2      , 4'd15     , 4'd3      , 4'd12     , 4'd14     , 4'd5      , 4'd11     , 4'd3      , 4'd8      , 4'd6      , 4'd4      , 4'd6      , 4'd12     , 4'd3      , 4'd6      , 4'd2      , 4'd12     , 4'd12     , 4'd6      , 4'd5      , 4'd11     , 4'd5      , 4'd13     , 4'd9      , 4'd4      , 4'd6      , 4'd13     , 4'd5      , 4'd11     , 4'd15     , 4'd1      , 4'd3      , 4'd13     , 4'd3      , 4'd10     , 4'd8      , 4'd14     , 4'd9      , 4'd5      , 4'd13     , 4'd5      , 4'd6      , 4'd0      , 4'd9      , 4'd14     , 4'd7       },
    '{ 4'd5      , 4'd15     , 4'd1      , 4'd5      , 4'd6      , 4'd12     , 4'd10     , 4'd10     , 4'd11     , 4'd6      , 4'd14     , 4'd14     , 4'd8      , 4'd7      , 4'd13     , 4'd5      , 4'd15     , 4'd11     , 4'd10     , 4'd3      , 4'd10     , 4'd2      , 4'd9      , 4'd11     , 4'd9      , 4'd3      , 4'd13     , 4'd14     , 4'd2      , 4'd5      , 4'd10     , 4'd4      , 4'd1      , 4'd5      , 4'd15     , 4'd14     , 4'd8      , 4'd3      , 4'd5      , 4'd8      , 4'd4      , 4'd10     , 4'd1      , 4'd7      , 4'd8      , 4'd1      , 4'd2      , 4'd1      , 4'd14     , 4'd1       },
    '{ 4'd7      , 4'd5      , 4'd11     , 4'd14     , 4'd0      , 4'd4      , 4'd15     , 4'd1      , 4'd1      , 4'd13     , 4'd12     , 4'd6      , 4'd14     , 4'd6      , 4'd0      , 4'd2      , 4'd3      , 4'd7      , 4'd12     , 4'd9      , 4'd14     , 4'd2      , 4'd11     , 4'd4      , 4'd9      , 4'd14     , 4'd0      , 4'd12     , 4'd6      , 4'd9      , 4'd2      , 4'd4      , 4'd7      , 4'd3      , 4'd0      , 4'd12     , 4'd5      , 4'd4      , 4'd13     , 4'd0      , 4'd13     , 4'd2      , 4'd3      , 4'd1      , 4'd7      , 4'd10     , 4'd1      , 4'd14     , 4'd13     , 4'd3       },
    '{ 4'd10     , 4'd4      , 4'd10     , 4'd1      , 4'd7      , 4'd4      , 4'd0      , 4'd10     , 4'd2      , 4'd12     , 4'd10     , 4'd7      , 4'd4      , 4'd0      , 4'd2      , 4'd6      , 4'd9      , 4'd2      , 4'd4      , 4'd12     , 4'd9      , 4'd9      , 4'd12     , 4'd5      , 4'd4      , 4'd10     , 4'd4      , 4'd9      , 4'd10     , 4'd12     , 4'd8      , 4'd1      , 4'd5      , 4'd7      , 4'd0      , 4'd10     , 4'd1      , 4'd10     , 4'd3      , 4'd9      , 4'd2      , 4'd8      , 4'd2      , 4'd4      , 4'd14     , 4'd12     , 4'd8      , 4'd2      , 4'd9      , 4'd8       }
  };

  assign weights_n2 = '{
    4'd7 ,
    4'd10,
    4'd11,
    4'd12,
    4'd8 ,
    4'd2 ,
    4'd3 ,
    4'd12,
    4'd3 ,
    4'd13,
    4'd6 
  };

  assign tanh = '{
    16'd16384,
    16'd59530,
    16'd53955,
    16'd63366,
    16'd38619,
    16'd46947,
    16'd43449,
    16'd61382,
    16'd52115,
    16'd58530,
    16'd2098,
    16'd47346,
    16'd37734,
    16'd2068,
    16'd6827,
    16'd12918
  };
endmodule
